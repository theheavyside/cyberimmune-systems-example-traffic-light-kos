component traffic_light.CStatus

endpoints {
    /* Declaration of a named implementation of the "Mode" interface. */
    mode : traffic_light.IStatus
}
